module Floating_point_unit(
    input clk,
    input wire [1:0] operation,
    input wire [15:0] op1,
    input wire [15:0] op2
);



endmodule